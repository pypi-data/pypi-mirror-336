/* Simple Top Module */
module simplemodule(
	input wire clk,
 	input wire reset	
    );
	   
endmodule

